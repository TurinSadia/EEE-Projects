-----------UVM Files------------ 

import uvm_pkg;
`include  uvm_macros.svh
`include params.sv
-----------RTL Files------------  
`include slave_rtl.sv
`include apb_rtl.sv
  
---------Customize Files--------
`include apb_interface.sv

`include apb_sequence_item.sv
`include apb_scoreboard.sv 

`include apb_sequencer.sv
`include apb_driver.sv
`include apb_monitor.sv
`include apb_agent.sv
`include apb_scoreboard.sv
`include apb_sequence.sv
`include apb_env.sv
`include apb_test.sv
`include apb_top.sv
